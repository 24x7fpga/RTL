`include "package.svh"
module $ARG (/*AUTOARG*/);
   // Outputs

   // Inputs


   /*AUTOREG*/
   /*AUTOWIRE*/

   <module> MOD1 (/*AUTOINST*/);

endmodule // $ARG
// Local Variables:
// Verilog-Library-Directories: (".")
// End:
