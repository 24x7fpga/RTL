`ifndef PACKAGE_SVH
 `define PACKAGE_SVH

// Define Timescale
 `timescale 1ns/1ns

// Define Clock
`define T 8  // 125MHz => Zybo Z7-20

`endif
