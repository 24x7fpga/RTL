`timescale 1ns/1ns
module spi_master #(parameter mode = 0) (/*AUTOARG*/);
   //outputs
   
endmodule // spi_master
// Local Variables: 
// Verilog-Library-Directories: (".")
// End:
