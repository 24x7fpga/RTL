`ifndef PACKAGE_SVH
 `define PACKAGE_SVH

// Define Timescale
 `timescale 1ns/1ns

// Define Clock
`define T     4'd8      // 125MHz => Zybo Z7-20
`define DVSR 12'd500    // 400kHz

`endif
