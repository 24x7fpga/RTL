kiran@Kirans-MacBook-Pro.local.2850